library verilog;
use verilog.vl_types.all;
entity shiftLeft226 is
    port(
        \in\            : in     vl_logic_vector(25 downto 0);
        \out\           : out    vl_logic_vector(27 downto 0)
    );
end shiftLeft226;
