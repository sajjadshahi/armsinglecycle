library verilog;
use verilog.vl_types.all;
entity testbranch is
end testbranch;
